`timescale 1ns / 1ps


module decoder4_16_tb;
reg a1,a2,a3,w,e;
wire [15:0]d;
decoder4_16 uut(a1,a2,a3,w,e,d);
initial
begin
#20 e=0; a1=0; a2=0; a3=0; w=0;
#40 e=1; a1=0; a2=0; a3=0; w=1;
#60 e=1; a1=0; a2=0; a3=1; w=0;
#80 e=1; a1=0; a2=0; a3=1; w=1;
#100 e=1; a1=0; a2=1; a3=0; w=0;
#120 e=1; a1=0; a2=1; a3=0; w=1;
#140 e=1; a1=0; a2=1; a3=1; w=0;
#160 e=1; a1=0; a2=1; a3=1; w=1;
#200 e=0; a1=1; a2=0; a3=0; w=1;
#220 e=0; a1=1; a2=0; a3=1; w=0;
#240 e=0; a1=1; a2=0; a3=1; w=1;
#260 e=0; a1=1; a2=1; a3=0; w=0;
#280 e=0; a1=1; a2=1; a3=0; w=1;
#300 e=0; a1=1; a2=1; a3=1; w=0;
#320 e=0; a1=1; a2=1; a3=1; w=1;


end
endmodule
